// Custom Module

 module rw_top();
 		

                 


	

endmodule
